    Mac OS X            	   2  ]     �                                      ATTR      �   �   �                  �   �  com.apple.acl.text     <   S  com.dropbox.attributes   !#acl 1
user:FFFFEEEE-DDDD-CCCC-BBBB-AAAA00000059:_spotlight:89:allow,inherited:read,execute,readattr,readextattr,readsecurity
 x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK����ʨ`�����(/���L#� ��r[[���Z �Q�